// FPGA Top Level

`default_nettype none

module top (
  // I/O ports
  input  logic hz100, reset,
  input  logic [20:0] pb,
  output logic [7:0] left, right,
         ss7, ss6, ss5, ss4, ss3, ss2, ss1, ss0,
  output logic red, green, blue,

  // UART ports
  output logic [7:0] txdata,
  input  logic [7:0] rxdata,
  output logic txclk, rxclk,
  input  logic txready, rxready
);
logic [31:0] out;
pc testpc(.clk(hz100), .nRST(~pb[19]), .ALUneg(1), .Zero(1), .iready(1), .PCaddr(out), .cuOP(6'b0), .rs1Read(32'b0), .signExtend(32'b0));
endmodule

