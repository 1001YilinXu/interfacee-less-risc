module request ();
    input logic CLK, nRST, 
    input logic [31:0] imemaddr, dmmaddr, dmmstore,
    input cuOPType cuOP;
endmodule